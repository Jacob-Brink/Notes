library verilog;
use verilog.vl_types.all;
entity Lab4BABY_vlg_vec_tst is
end Lab4BABY_vlg_vec_tst;
