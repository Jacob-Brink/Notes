library verilog;
use verilog.vl_types.all;
entity Lab4BABY_vlg_check_tst is
    port(
        Unit0LED        : in     vl_logic;
        Unit1LED        : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab4BABY_vlg_check_tst;
