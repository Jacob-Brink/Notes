library verilog;
use verilog.vl_types.all;
entity Lab2_SectionB_vlg_check_tst is
    port(
        D               : in     vl_logic;
        SimpD           : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end Lab2_SectionB_vlg_check_tst;
