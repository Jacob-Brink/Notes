library verilog;
use verilog.vl_types.all;
entity Lab3_vlg_vec_tst is
end Lab3_vlg_vec_tst;
